magic
tech scmos
timestamp 1703850560
<< nwell >>
rect 175 -92 448 -67
<< ntransistor >>
rect 186 -123 188 -119
rect 204 -123 206 -119
rect 222 -123 224 -119
rect 238 -123 240 -119
rect 254 -123 256 -119
rect 275 -123 277 -119
rect 293 -123 295 -119
rect 311 -123 313 -119
rect 327 -123 329 -119
rect 343 -123 345 -119
rect 367 -123 369 -119
rect 385 -123 387 -119
rect 403 -123 405 -119
rect 419 -123 421 -119
rect 435 -123 437 -119
<< ptransistor >>
rect 186 -86 188 -78
rect 204 -86 206 -78
rect 222 -86 224 -78
rect 238 -86 240 -78
rect 254 -86 256 -78
rect 275 -86 277 -78
rect 293 -86 295 -78
rect 311 -86 313 -78
rect 327 -86 329 -78
rect 343 -86 345 -78
rect 367 -86 369 -78
rect 385 -86 387 -78
rect 403 -86 405 -78
rect 419 -86 421 -78
rect 435 -86 437 -78
<< ndiffusion >>
rect 185 -123 186 -119
rect 188 -123 189 -119
rect 203 -123 204 -119
rect 206 -123 207 -119
rect 221 -123 222 -119
rect 224 -123 225 -119
rect 237 -123 238 -119
rect 240 -123 241 -119
rect 253 -123 254 -119
rect 256 -123 257 -119
rect 274 -123 275 -119
rect 277 -123 278 -119
rect 292 -123 293 -119
rect 295 -123 296 -119
rect 310 -123 311 -119
rect 313 -123 314 -119
rect 326 -123 327 -119
rect 329 -123 330 -119
rect 342 -123 343 -119
rect 345 -123 346 -119
rect 366 -123 367 -119
rect 369 -123 370 -119
rect 384 -123 385 -119
rect 387 -123 388 -119
rect 402 -123 403 -119
rect 405 -123 406 -119
rect 418 -123 419 -119
rect 421 -123 422 -119
rect 434 -123 435 -119
rect 437 -123 438 -119
<< pdiffusion >>
rect 185 -86 186 -78
rect 188 -86 189 -78
rect 203 -86 204 -78
rect 206 -86 207 -78
rect 221 -86 222 -78
rect 224 -86 225 -78
rect 237 -86 238 -78
rect 240 -86 241 -78
rect 253 -86 254 -78
rect 256 -86 257 -78
rect 274 -86 275 -78
rect 277 -86 278 -78
rect 292 -86 293 -78
rect 295 -86 296 -78
rect 310 -86 311 -78
rect 313 -86 314 -78
rect 326 -86 327 -78
rect 329 -86 330 -78
rect 342 -86 343 -78
rect 345 -86 346 -78
rect 366 -86 367 -78
rect 369 -86 370 -78
rect 384 -86 385 -78
rect 387 -86 388 -78
rect 402 -86 403 -78
rect 405 -86 406 -78
rect 418 -86 419 -78
rect 421 -86 422 -78
rect 434 -86 435 -78
rect 437 -86 438 -78
<< ndcontact >>
rect 181 -123 185 -119
rect 189 -123 193 -119
rect 199 -123 203 -119
rect 207 -123 211 -119
rect 217 -123 221 -119
rect 225 -123 229 -119
rect 233 -123 237 -119
rect 241 -123 245 -119
rect 249 -123 253 -119
rect 257 -123 261 -119
rect 270 -123 274 -119
rect 278 -123 282 -119
rect 288 -123 292 -119
rect 296 -123 300 -119
rect 306 -123 310 -119
rect 314 -123 318 -119
rect 322 -123 326 -119
rect 330 -123 334 -119
rect 338 -123 342 -119
rect 346 -123 350 -119
rect 362 -123 366 -119
rect 370 -123 374 -119
rect 380 -123 384 -119
rect 388 -123 392 -119
rect 398 -123 402 -119
rect 406 -123 410 -119
rect 414 -123 418 -119
rect 422 -123 426 -119
rect 430 -123 434 -119
rect 438 -123 442 -119
<< pdcontact >>
rect 181 -86 185 -78
rect 189 -86 193 -78
rect 199 -86 203 -78
rect 207 -86 211 -78
rect 217 -86 221 -78
rect 225 -86 229 -78
rect 233 -86 237 -78
rect 241 -86 245 -78
rect 249 -86 253 -78
rect 257 -86 261 -78
rect 270 -86 274 -78
rect 278 -86 282 -78
rect 288 -86 292 -78
rect 296 -86 300 -78
rect 306 -86 310 -78
rect 314 -86 318 -78
rect 322 -86 326 -78
rect 330 -86 334 -78
rect 338 -86 342 -78
rect 346 -86 350 -78
rect 362 -86 366 -78
rect 370 -86 374 -78
rect 380 -86 384 -78
rect 388 -86 392 -78
rect 398 -86 402 -78
rect 406 -86 410 -78
rect 414 -86 418 -78
rect 422 -86 426 -78
rect 430 -86 434 -78
rect 438 -86 442 -78
<< polysilicon >>
rect 186 -78 188 -75
rect 204 -78 206 -75
rect 222 -78 224 -75
rect 238 -78 240 -75
rect 254 -78 256 -75
rect 275 -78 277 -75
rect 293 -78 295 -75
rect 311 -78 313 -75
rect 327 -78 329 -75
rect 343 -78 345 -75
rect 367 -78 369 -75
rect 385 -78 387 -75
rect 403 -78 405 -75
rect 419 -78 421 -75
rect 435 -78 437 -75
rect 186 -119 188 -86
rect 204 -119 206 -86
rect 222 -119 224 -86
rect 238 -119 240 -86
rect 254 -119 256 -86
rect 275 -119 277 -86
rect 293 -119 295 -86
rect 311 -119 313 -86
rect 327 -119 329 -86
rect 343 -119 345 -86
rect 367 -119 369 -86
rect 385 -119 387 -86
rect 403 -119 405 -86
rect 419 -119 421 -86
rect 435 -119 437 -86
rect 186 -126 188 -123
rect 204 -126 206 -123
rect 222 -126 224 -123
rect 238 -126 240 -123
rect 254 -126 256 -123
rect 275 -126 277 -123
rect 293 -126 295 -123
rect 311 -126 313 -123
rect 327 -126 329 -123
rect 343 -126 345 -123
rect 367 -126 369 -123
rect 385 -126 387 -123
rect 403 -126 405 -123
rect 419 -126 421 -123
rect 435 -126 437 -123
<< polycontact >>
rect 200 -100 204 -96
rect 188 -109 192 -105
rect 218 -100 222 -96
rect 240 -109 244 -105
rect 256 -105 260 -101
rect 289 -100 293 -96
rect 277 -109 281 -105
rect 307 -98 311 -94
rect 329 -109 333 -105
rect 345 -105 349 -101
rect 381 -100 385 -96
rect 369 -109 373 -105
rect 399 -98 403 -94
rect 421 -109 425 -105
rect 437 -105 441 -101
<< metal1 >>
rect 176 -74 446 -69
rect 181 -78 185 -74
rect 199 -78 203 -74
rect 257 -78 261 -74
rect 211 -80 217 -78
rect 211 -85 212 -80
rect 211 -86 217 -85
rect 189 -89 193 -86
rect 207 -89 211 -86
rect 189 -93 211 -89
rect 185 -100 200 -96
rect 225 -97 229 -86
rect 241 -97 245 -86
rect 225 -101 245 -97
rect 270 -78 274 -74
rect 288 -78 292 -74
rect 346 -78 350 -74
rect 300 -80 306 -78
rect 300 -85 301 -80
rect 300 -86 306 -85
rect 225 -112 229 -101
rect 249 -105 253 -86
rect 278 -89 282 -86
rect 296 -89 300 -86
rect 278 -93 300 -89
rect 256 -101 260 -96
rect 285 -100 289 -96
rect 303 -98 307 -94
rect 314 -97 318 -86
rect 330 -97 334 -86
rect 314 -101 334 -97
rect 362 -78 366 -74
rect 380 -78 384 -74
rect 438 -78 442 -74
rect 392 -80 398 -78
rect 392 -85 393 -80
rect 392 -86 398 -85
rect 244 -109 253 -105
rect 176 -116 245 -112
rect 181 -119 185 -116
rect 241 -119 245 -116
rect 193 -123 199 -119
rect 207 -127 211 -123
rect 229 -123 233 -119
rect 249 -119 253 -109
rect 314 -112 318 -101
rect 338 -105 342 -86
rect 370 -89 374 -86
rect 388 -89 392 -86
rect 370 -93 392 -89
rect 377 -100 381 -96
rect 395 -98 399 -94
rect 406 -97 410 -86
rect 422 -97 426 -86
rect 406 -101 426 -97
rect 333 -109 342 -105
rect 274 -116 334 -112
rect 270 -119 274 -117
rect 330 -119 334 -116
rect 282 -123 288 -119
rect 217 -127 221 -123
rect 257 -127 261 -123
rect 296 -127 300 -123
rect 318 -123 322 -119
rect 338 -119 342 -109
rect 406 -112 410 -101
rect 430 -105 434 -86
rect 437 -101 441 -96
rect 425 -109 434 -105
rect 357 -117 358 -112
rect 363 -116 426 -112
rect 363 -117 366 -116
rect 362 -119 366 -117
rect 422 -119 426 -116
rect 374 -123 380 -119
rect 306 -127 310 -123
rect 346 -127 350 -123
rect 388 -127 392 -123
rect 410 -123 414 -119
rect 430 -119 434 -109
rect 398 -127 402 -123
rect 438 -127 442 -123
rect 176 -132 444 -127
<< m2contact >>
rect 212 -85 217 -80
rect 180 -101 185 -96
rect 213 -101 218 -96
rect 232 -91 237 -86
rect 301 -85 306 -80
rect 192 -109 197 -104
rect 321 -91 326 -86
rect 393 -85 398 -80
rect 260 -106 265 -101
rect 281 -109 286 -104
rect 413 -91 418 -86
rect 349 -106 354 -101
rect 373 -109 378 -104
rect 269 -117 274 -112
rect 441 -106 446 -101
rect 358 -117 363 -112
<< metal2 >>
rect 203 -75 362 -71
rect 203 -96 207 -75
rect 212 -86 217 -85
rect 301 -86 306 -85
rect 212 -91 232 -86
rect 301 -91 321 -86
rect 203 -100 213 -96
rect 180 -113 185 -101
rect 197 -106 260 -105
rect 197 -109 265 -106
rect 286 -106 349 -105
rect 286 -109 354 -106
rect 180 -117 269 -113
rect 350 -127 354 -109
rect 358 -112 362 -75
rect 393 -86 398 -85
rect 393 -91 413 -86
rect 378 -106 441 -105
rect 378 -109 446 -106
rect 442 -127 446 -109
rect 350 -131 446 -127
<< labels >>
rlabel metal1 273 -130 273 -130 1 Gnd
rlabel metal1 275 -71 275 -71 1 Vdd
rlabel metal1 395 -98 395 -94 1 D0
rlabel metal1 365 -130 365 -130 1 Gnd
rlabel metal1 367 -71 367 -71 1 Vdd
rlabel metal1 176 -116 176 -112 3 Y
rlabel metal1 184 -130 184 -130 1 Gnd
rlabel metal1 186 -71 186 -71 1 Vdd
rlabel metal1 256 -96 260 -96 1 S1
rlabel metal1 437 -96 441 -96 1 S0
rlabel metal1 285 -100 285 -96 1 D3
rlabel metal1 303 -98 303 -94 1 D1
rlabel metal1 377 -100 377 -96 1 D2
<< end >>
