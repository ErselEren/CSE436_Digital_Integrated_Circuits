magic
tech scmos
timestamp 1702654670
<< nwell >>
rect -38 263 562 288
rect -38 196 563 221
rect -38 129 563 154
rect -38 62 563 87
<< ntransistor >>
rect -27 232 -25 236
rect -1 232 1 236
rect 11 232 13 236
rect 31 232 33 236
rect 57 232 59 236
rect 83 232 85 236
rect 95 232 97 236
rect 115 232 117 236
rect 134 232 136 236
rect 145 232 147 236
rect 165 232 167 236
rect 185 232 187 236
rect 195 232 197 236
rect 215 232 217 236
rect 250 232 252 236
rect 276 232 278 236
rect 288 232 290 236
rect 308 232 310 236
rect 334 232 336 236
rect 360 232 362 236
rect 372 232 374 236
rect 392 232 394 236
rect 411 232 413 236
rect 422 232 424 236
rect 442 232 444 236
rect 462 232 464 236
rect 472 232 474 236
rect 492 232 494 236
rect 517 232 519 236
rect 528 232 530 236
rect 548 232 550 236
rect -27 165 -25 169
rect -1 165 1 169
rect 11 165 13 169
rect 31 165 33 169
rect 57 165 59 169
rect 83 165 85 169
rect 95 165 97 169
rect 115 165 117 169
rect 134 165 136 169
rect 145 165 147 169
rect 165 165 167 169
rect 185 165 187 169
rect 195 165 197 169
rect 215 165 217 169
rect 250 165 252 169
rect 276 165 278 169
rect 288 165 290 169
rect 308 165 310 169
rect 334 165 336 169
rect 360 165 362 169
rect 372 165 374 169
rect 392 165 394 169
rect 411 165 413 169
rect 422 165 424 169
rect 442 165 444 169
rect 462 165 464 169
rect 472 165 474 169
rect 492 165 494 169
rect 517 165 519 169
rect 528 165 530 169
rect 548 165 550 169
rect -27 98 -25 102
rect -1 98 1 102
rect 11 98 13 102
rect 31 98 33 102
rect 57 98 59 102
rect 83 98 85 102
rect 95 98 97 102
rect 115 98 117 102
rect 134 98 136 102
rect 145 98 147 102
rect 165 98 167 102
rect 185 98 187 102
rect 195 98 197 102
rect 215 98 217 102
rect 250 98 252 102
rect 276 98 278 102
rect 288 98 290 102
rect 308 98 310 102
rect 334 98 336 102
rect 360 98 362 102
rect 372 98 374 102
rect 392 98 394 102
rect 411 98 413 102
rect 422 98 424 102
rect 442 98 444 102
rect 462 98 464 102
rect 472 98 474 102
rect 492 98 494 102
rect 517 98 519 102
rect 528 98 530 102
rect 548 98 550 102
rect -27 31 -25 35
rect -1 31 1 35
rect 11 31 13 35
rect 31 31 33 35
rect 57 31 59 35
rect 83 31 85 35
rect 95 31 97 35
rect 115 31 117 35
rect 134 31 136 35
rect 145 31 147 35
rect 165 31 167 35
rect 185 31 187 35
rect 195 31 197 35
rect 215 31 217 35
rect 250 31 252 35
rect 276 31 278 35
rect 288 31 290 35
rect 308 31 310 35
rect 334 31 336 35
rect 360 31 362 35
rect 372 31 374 35
rect 392 31 394 35
rect 411 31 413 35
rect 422 31 424 35
rect 442 31 444 35
rect 462 31 464 35
rect 472 31 474 35
rect 492 31 494 35
rect 517 31 519 35
rect 528 31 530 35
rect 548 31 550 35
<< ptransistor >>
rect -27 269 -25 277
rect -1 269 1 277
rect 11 269 13 277
rect 31 269 33 277
rect 57 269 59 277
rect 83 269 85 277
rect 95 269 97 277
rect 115 269 117 277
rect 134 269 136 277
rect 145 269 147 277
rect 165 269 167 277
rect 185 269 187 277
rect 195 269 197 277
rect 215 269 217 277
rect 250 269 252 277
rect 276 269 278 277
rect 288 269 290 277
rect 308 269 310 277
rect 334 269 336 277
rect 360 269 362 277
rect 372 269 374 277
rect 392 269 394 277
rect 411 269 413 277
rect 422 269 424 277
rect 442 269 444 277
rect 462 269 464 277
rect 472 269 474 277
rect 492 269 494 277
rect 517 269 519 277
rect 528 269 530 277
rect 548 269 550 277
rect -27 202 -25 210
rect -1 202 1 210
rect 11 202 13 210
rect 31 202 33 210
rect 57 202 59 210
rect 83 202 85 210
rect 95 202 97 210
rect 115 202 117 210
rect 134 202 136 210
rect 145 202 147 210
rect 165 202 167 210
rect 185 202 187 210
rect 195 202 197 210
rect 215 202 217 210
rect 250 202 252 210
rect 276 202 278 210
rect 288 202 290 210
rect 308 202 310 210
rect 334 202 336 210
rect 360 202 362 210
rect 372 202 374 210
rect 392 202 394 210
rect 411 202 413 210
rect 422 202 424 210
rect 442 202 444 210
rect 462 202 464 210
rect 472 202 474 210
rect 492 202 494 210
rect 517 202 519 210
rect 528 202 530 210
rect 548 202 550 210
rect -27 135 -25 143
rect -1 135 1 143
rect 11 135 13 143
rect 31 135 33 143
rect 57 135 59 143
rect 83 135 85 143
rect 95 135 97 143
rect 115 135 117 143
rect 134 135 136 143
rect 145 135 147 143
rect 165 135 167 143
rect 185 135 187 143
rect 195 135 197 143
rect 215 135 217 143
rect 250 135 252 143
rect 276 135 278 143
rect 288 135 290 143
rect 308 135 310 143
rect 334 135 336 143
rect 360 135 362 143
rect 372 135 374 143
rect 392 135 394 143
rect 411 135 413 143
rect 422 135 424 143
rect 442 135 444 143
rect 462 135 464 143
rect 472 135 474 143
rect 492 135 494 143
rect 517 135 519 143
rect 528 135 530 143
rect 548 135 550 143
rect -27 68 -25 76
rect -1 68 1 76
rect 11 68 13 76
rect 31 68 33 76
rect 57 68 59 76
rect 83 68 85 76
rect 95 68 97 76
rect 115 68 117 76
rect 134 68 136 76
rect 145 68 147 76
rect 165 68 167 76
rect 185 68 187 76
rect 195 68 197 76
rect 215 68 217 76
rect 250 68 252 76
rect 276 68 278 76
rect 288 68 290 76
rect 308 68 310 76
rect 334 68 336 76
rect 360 68 362 76
rect 372 68 374 76
rect 392 68 394 76
rect 411 68 413 76
rect 422 68 424 76
rect 442 68 444 76
rect 462 68 464 76
rect 472 68 474 76
rect 492 68 494 76
rect 517 68 519 76
rect 528 68 530 76
rect 548 68 550 76
<< ndiffusion >>
rect -28 232 -27 236
rect -25 232 -24 236
rect -2 232 -1 236
rect 1 232 11 236
rect 13 232 14 236
rect 30 232 31 236
rect 33 232 34 236
rect 56 232 57 236
rect 59 232 60 236
rect 82 232 83 236
rect 85 232 95 236
rect 97 232 98 236
rect 114 232 115 236
rect 117 232 118 236
rect 133 232 134 236
rect 136 232 140 236
rect 144 232 145 236
rect 147 232 148 236
rect 164 232 165 236
rect 167 232 168 236
rect 184 232 185 236
rect 187 232 195 236
rect 197 232 198 236
rect 214 232 215 236
rect 217 232 218 236
rect 249 232 250 236
rect 252 232 253 236
rect 275 232 276 236
rect 278 232 288 236
rect 290 232 291 236
rect 307 232 308 236
rect 310 232 311 236
rect 333 232 334 236
rect 336 232 337 236
rect 359 232 360 236
rect 362 232 372 236
rect 374 232 375 236
rect 391 232 392 236
rect 394 232 395 236
rect 410 232 411 236
rect 413 232 417 236
rect 421 232 422 236
rect 424 232 425 236
rect 441 232 442 236
rect 444 232 445 236
rect 461 232 462 236
rect 464 232 472 236
rect 474 232 475 236
rect 491 232 492 236
rect 494 232 495 236
rect 516 232 517 236
rect 519 232 523 236
rect 527 232 528 236
rect 530 232 531 236
rect 547 232 548 236
rect 550 232 551 236
rect -28 165 -27 169
rect -25 165 -24 169
rect -2 165 -1 169
rect 1 165 11 169
rect 13 165 14 169
rect 30 165 31 169
rect 33 165 34 169
rect 56 165 57 169
rect 59 165 60 169
rect 82 165 83 169
rect 85 165 95 169
rect 97 165 98 169
rect 114 165 115 169
rect 117 165 118 169
rect 133 165 134 169
rect 136 165 140 169
rect 144 165 145 169
rect 147 165 148 169
rect 164 165 165 169
rect 167 165 168 169
rect 184 165 185 169
rect 187 165 195 169
rect 197 165 198 169
rect 214 165 215 169
rect 217 165 218 169
rect 249 165 250 169
rect 252 165 253 169
rect 275 165 276 169
rect 278 165 288 169
rect 290 165 291 169
rect 307 165 308 169
rect 310 165 311 169
rect 333 165 334 169
rect 336 165 337 169
rect 359 165 360 169
rect 362 165 372 169
rect 374 165 375 169
rect 391 165 392 169
rect 394 165 395 169
rect 410 165 411 169
rect 413 165 417 169
rect 421 165 422 169
rect 424 165 425 169
rect 441 165 442 169
rect 444 165 445 169
rect 461 165 462 169
rect 464 165 472 169
rect 474 165 475 169
rect 491 165 492 169
rect 494 165 495 169
rect 516 165 517 169
rect 519 165 523 169
rect 527 165 528 169
rect 530 165 531 169
rect 547 165 548 169
rect 550 165 551 169
rect -28 98 -27 102
rect -25 98 -24 102
rect -2 98 -1 102
rect 1 98 11 102
rect 13 98 14 102
rect 30 98 31 102
rect 33 98 34 102
rect 56 98 57 102
rect 59 98 60 102
rect 82 98 83 102
rect 85 98 95 102
rect 97 98 98 102
rect 114 98 115 102
rect 117 98 118 102
rect 133 98 134 102
rect 136 98 140 102
rect 144 98 145 102
rect 147 98 148 102
rect 164 98 165 102
rect 167 98 168 102
rect 184 98 185 102
rect 187 98 195 102
rect 197 98 198 102
rect 214 98 215 102
rect 217 98 218 102
rect 249 98 250 102
rect 252 98 253 102
rect 275 98 276 102
rect 278 98 288 102
rect 290 98 291 102
rect 307 98 308 102
rect 310 98 311 102
rect 333 98 334 102
rect 336 98 337 102
rect 359 98 360 102
rect 362 98 372 102
rect 374 98 375 102
rect 391 98 392 102
rect 394 98 395 102
rect 410 98 411 102
rect 413 98 417 102
rect 421 98 422 102
rect 424 98 425 102
rect 441 98 442 102
rect 444 98 445 102
rect 461 98 462 102
rect 464 98 472 102
rect 474 98 475 102
rect 491 98 492 102
rect 494 98 495 102
rect 516 98 517 102
rect 519 98 523 102
rect 527 98 528 102
rect 530 98 531 102
rect 547 98 548 102
rect 550 98 551 102
rect -28 31 -27 35
rect -25 31 -24 35
rect -2 31 -1 35
rect 1 31 11 35
rect 13 31 14 35
rect 30 31 31 35
rect 33 31 34 35
rect 56 31 57 35
rect 59 31 60 35
rect 82 31 83 35
rect 85 31 95 35
rect 97 31 98 35
rect 114 31 115 35
rect 117 31 118 35
rect 133 31 134 35
rect 136 31 140 35
rect 144 31 145 35
rect 147 31 148 35
rect 164 31 165 35
rect 167 31 168 35
rect 184 31 185 35
rect 187 31 195 35
rect 197 31 198 35
rect 214 31 215 35
rect 217 31 218 35
rect 249 31 250 35
rect 252 31 253 35
rect 275 31 276 35
rect 278 31 288 35
rect 290 31 291 35
rect 307 31 308 35
rect 310 31 311 35
rect 333 31 334 35
rect 336 31 337 35
rect 359 31 360 35
rect 362 31 372 35
rect 374 31 375 35
rect 391 31 392 35
rect 394 31 395 35
rect 410 31 411 35
rect 413 31 417 35
rect 421 31 422 35
rect 424 31 425 35
rect 441 31 442 35
rect 444 31 445 35
rect 461 31 462 35
rect 464 31 472 35
rect 474 31 475 35
rect 491 31 492 35
rect 494 31 495 35
rect 516 31 517 35
rect 519 31 523 35
rect 527 31 528 35
rect 530 31 531 35
rect 547 31 548 35
rect 550 31 551 35
<< pdiffusion >>
rect -28 269 -27 277
rect -25 269 -24 277
rect -20 269 -18 277
rect -2 269 -1 277
rect 1 269 2 277
rect 6 269 11 277
rect 13 269 14 277
rect 30 269 31 277
rect 33 269 34 277
rect 38 269 40 277
rect 56 269 57 277
rect 59 269 60 277
rect 64 269 66 277
rect 82 269 83 277
rect 85 269 86 277
rect 90 269 95 277
rect 97 269 98 277
rect 114 269 115 277
rect 117 269 118 277
rect 122 269 124 277
rect 133 269 134 277
rect 136 269 145 277
rect 147 269 148 277
rect 164 269 165 277
rect 167 269 168 277
rect 172 269 174 277
rect 184 269 185 277
rect 187 269 188 277
rect 194 269 195 277
rect 197 269 198 277
rect 214 269 215 277
rect 217 269 218 277
rect 222 269 224 277
rect 249 269 250 277
rect 252 269 253 277
rect 257 269 259 277
rect 275 269 276 277
rect 278 269 279 277
rect 283 269 288 277
rect 290 269 291 277
rect 307 269 308 277
rect 310 269 311 277
rect 315 269 317 277
rect 333 269 334 277
rect 336 269 337 277
rect 341 269 343 277
rect 359 269 360 277
rect 362 269 363 277
rect 367 269 372 277
rect 374 269 375 277
rect 391 269 392 277
rect 394 269 395 277
rect 399 269 401 277
rect 410 269 411 277
rect 413 269 422 277
rect 424 269 425 277
rect 441 269 442 277
rect 444 269 445 277
rect 449 269 451 277
rect 461 269 462 277
rect 464 269 465 277
rect 471 269 472 277
rect 474 269 475 277
rect 491 269 492 277
rect 494 269 495 277
rect 499 269 501 277
rect 516 269 517 277
rect 519 269 528 277
rect 530 269 531 277
rect 547 269 548 277
rect 550 269 551 277
rect 555 269 556 277
rect -28 202 -27 210
rect -25 202 -24 210
rect -20 202 -18 210
rect -2 202 -1 210
rect 1 202 2 210
rect 6 202 11 210
rect 13 202 14 210
rect 30 202 31 210
rect 33 202 34 210
rect 38 202 40 210
rect 56 202 57 210
rect 59 202 60 210
rect 64 202 66 210
rect 82 202 83 210
rect 85 202 86 210
rect 90 202 95 210
rect 97 202 98 210
rect 114 202 115 210
rect 117 202 118 210
rect 122 202 124 210
rect 133 202 134 210
rect 136 202 145 210
rect 147 202 148 210
rect 164 202 165 210
rect 167 202 168 210
rect 172 202 174 210
rect 184 202 185 210
rect 187 202 188 210
rect 194 202 195 210
rect 197 202 198 210
rect 214 202 215 210
rect 217 202 218 210
rect 222 202 224 210
rect 249 202 250 210
rect 252 202 253 210
rect 257 202 259 210
rect 275 202 276 210
rect 278 202 279 210
rect 283 202 288 210
rect 290 202 291 210
rect 307 202 308 210
rect 310 202 311 210
rect 315 202 317 210
rect 333 202 334 210
rect 336 202 337 210
rect 341 202 343 210
rect 359 202 360 210
rect 362 202 363 210
rect 367 202 372 210
rect 374 202 375 210
rect 391 202 392 210
rect 394 202 395 210
rect 399 202 401 210
rect 410 202 411 210
rect 413 202 422 210
rect 424 202 425 210
rect 441 202 442 210
rect 444 202 445 210
rect 449 202 451 210
rect 461 202 462 210
rect 464 202 465 210
rect 471 202 472 210
rect 474 202 475 210
rect 491 202 492 210
rect 494 202 495 210
rect 499 202 501 210
rect 516 202 517 210
rect 519 202 528 210
rect 530 202 531 210
rect 547 202 548 210
rect 550 202 551 210
rect 555 202 557 210
rect -28 135 -27 143
rect -25 135 -24 143
rect -20 135 -18 143
rect -2 135 -1 143
rect 1 135 2 143
rect 6 135 11 143
rect 13 135 14 143
rect 30 135 31 143
rect 33 135 34 143
rect 38 135 40 143
rect 56 135 57 143
rect 59 135 60 143
rect 64 135 66 143
rect 82 135 83 143
rect 85 135 86 143
rect 90 135 95 143
rect 97 135 98 143
rect 114 135 115 143
rect 117 135 118 143
rect 122 135 124 143
rect 133 135 134 143
rect 136 135 145 143
rect 147 135 148 143
rect 164 135 165 143
rect 167 135 168 143
rect 172 135 174 143
rect 184 135 185 143
rect 187 135 188 143
rect 194 135 195 143
rect 197 135 198 143
rect 214 135 215 143
rect 217 135 218 143
rect 222 135 224 143
rect 249 135 250 143
rect 252 135 253 143
rect 257 135 259 143
rect 275 135 276 143
rect 278 135 279 143
rect 283 135 288 143
rect 290 135 291 143
rect 307 135 308 143
rect 310 135 311 143
rect 315 135 317 143
rect 333 135 334 143
rect 336 135 337 143
rect 341 135 343 143
rect 359 135 360 143
rect 362 135 363 143
rect 367 135 372 143
rect 374 135 375 143
rect 391 135 392 143
rect 394 135 395 143
rect 399 135 401 143
rect 410 135 411 143
rect 413 135 422 143
rect 424 135 425 143
rect 441 135 442 143
rect 444 135 445 143
rect 449 135 451 143
rect 461 135 462 143
rect 464 135 465 143
rect 471 135 472 143
rect 474 135 475 143
rect 491 135 492 143
rect 494 135 495 143
rect 499 135 501 143
rect 516 135 517 143
rect 519 135 528 143
rect 530 135 531 143
rect 547 135 548 143
rect 550 135 551 143
rect 555 135 557 143
rect -28 68 -27 76
rect -25 68 -24 76
rect -20 68 -18 76
rect -2 68 -1 76
rect 1 68 2 76
rect 6 68 11 76
rect 13 68 14 76
rect 30 68 31 76
rect 33 68 34 76
rect 38 68 40 76
rect 56 68 57 76
rect 59 68 60 76
rect 64 68 66 76
rect 82 68 83 76
rect 85 68 86 76
rect 90 68 95 76
rect 97 68 98 76
rect 114 68 115 76
rect 117 68 118 76
rect 122 68 124 76
rect 133 68 134 76
rect 136 68 145 76
rect 147 68 148 76
rect 164 68 165 76
rect 167 68 168 76
rect 172 68 174 76
rect 184 68 185 76
rect 187 68 188 76
rect 194 68 195 76
rect 197 68 198 76
rect 214 68 215 76
rect 217 68 218 76
rect 222 68 224 76
rect 249 68 250 76
rect 252 68 253 76
rect 257 68 259 76
rect 275 68 276 76
rect 278 68 279 76
rect 283 68 288 76
rect 290 68 291 76
rect 307 68 308 76
rect 310 68 311 76
rect 315 68 317 76
rect 333 68 334 76
rect 336 68 337 76
rect 341 68 343 76
rect 359 68 360 76
rect 362 68 363 76
rect 367 68 372 76
rect 374 68 375 76
rect 391 68 392 76
rect 394 68 395 76
rect 399 68 401 76
rect 410 68 411 76
rect 413 68 422 76
rect 424 68 425 76
rect 441 68 442 76
rect 444 68 445 76
rect 449 68 451 76
rect 461 68 462 76
rect 464 68 465 76
rect 471 68 472 76
rect 474 68 475 76
rect 491 68 492 76
rect 494 68 495 76
rect 499 68 501 76
rect 516 68 517 76
rect 519 68 528 76
rect 530 68 531 76
rect 547 68 548 76
rect 550 68 551 76
rect 555 68 557 76
<< ndcontact >>
rect -32 232 -28 236
rect -24 232 -20 236
rect -6 232 -2 236
rect 14 232 18 236
rect 26 232 30 236
rect 34 232 38 236
rect 52 232 56 236
rect 60 232 64 236
rect 78 232 82 236
rect 98 232 102 236
rect 110 232 114 236
rect 118 232 122 236
rect 129 232 133 236
rect 140 232 144 236
rect 148 232 152 236
rect 160 232 164 236
rect 168 232 172 236
rect 180 232 184 236
rect 198 232 202 236
rect 210 232 214 236
rect 218 232 222 236
rect 245 232 249 236
rect 253 232 257 236
rect 271 232 275 236
rect 291 232 295 236
rect 303 232 307 236
rect 311 232 315 236
rect 329 232 333 236
rect 337 232 341 236
rect 355 232 359 236
rect 375 232 379 236
rect 387 232 391 236
rect 395 232 399 236
rect 406 232 410 236
rect 417 232 421 236
rect 425 232 429 236
rect 437 232 441 236
rect 445 232 449 236
rect 457 232 461 236
rect 475 232 479 236
rect 487 232 491 236
rect 495 232 499 236
rect 512 232 516 236
rect 523 232 527 236
rect 531 232 535 236
rect 543 232 547 236
rect 551 232 555 236
rect -32 165 -28 169
rect -24 165 -20 169
rect -6 165 -2 169
rect 14 165 18 169
rect 26 165 30 169
rect 34 165 38 169
rect 52 165 56 169
rect 60 165 64 169
rect 78 165 82 169
rect 98 165 102 169
rect 110 165 114 169
rect 118 165 122 169
rect 129 165 133 169
rect 140 165 144 169
rect 148 165 152 169
rect 160 165 164 169
rect 168 165 172 169
rect 180 165 184 169
rect 198 165 202 169
rect 210 165 214 169
rect 218 165 222 169
rect 245 165 249 169
rect 253 165 257 169
rect 271 165 275 169
rect 291 165 295 169
rect 303 165 307 169
rect 311 165 315 169
rect 329 165 333 169
rect 337 165 341 169
rect 355 165 359 169
rect 375 165 379 169
rect 387 165 391 169
rect 395 165 399 169
rect 406 165 410 169
rect 417 165 421 169
rect 425 165 429 169
rect 437 165 441 169
rect 445 165 449 169
rect 457 165 461 169
rect 475 165 479 169
rect 487 165 491 169
rect 495 165 499 169
rect 512 165 516 169
rect 523 165 527 169
rect 531 165 535 169
rect 543 165 547 169
rect 551 165 555 169
rect -32 98 -28 102
rect -24 98 -20 102
rect -6 98 -2 102
rect 14 98 18 102
rect 26 98 30 102
rect 34 98 38 102
rect 52 98 56 102
rect 60 98 64 102
rect 78 98 82 102
rect 98 98 102 102
rect 110 98 114 102
rect 118 98 122 102
rect 129 98 133 102
rect 140 98 144 102
rect 148 98 152 102
rect 160 98 164 102
rect 168 98 172 102
rect 180 98 184 102
rect 198 98 202 102
rect 210 98 214 102
rect 218 98 222 102
rect 245 98 249 102
rect 253 98 257 102
rect 271 98 275 102
rect 291 98 295 102
rect 303 98 307 102
rect 311 98 315 102
rect 329 98 333 102
rect 337 98 341 102
rect 355 98 359 102
rect 375 98 379 102
rect 387 98 391 102
rect 395 98 399 102
rect 406 98 410 102
rect 417 98 421 102
rect 425 98 429 102
rect 437 98 441 102
rect 445 98 449 102
rect 457 98 461 102
rect 475 98 479 102
rect 487 98 491 102
rect 495 98 499 102
rect 512 98 516 102
rect 523 98 527 102
rect 531 98 535 102
rect 543 98 547 102
rect 551 98 555 102
rect -32 31 -28 35
rect -24 31 -20 35
rect -6 31 -2 35
rect 14 31 18 35
rect 26 31 30 35
rect 34 31 38 35
rect 52 31 56 35
rect 60 31 64 35
rect 78 31 82 35
rect 98 31 102 35
rect 110 31 114 35
rect 118 31 122 35
rect 129 31 133 35
rect 140 31 144 35
rect 148 31 152 35
rect 160 31 164 35
rect 168 31 172 35
rect 180 31 184 35
rect 198 31 202 35
rect 210 31 214 35
rect 218 31 222 35
rect 245 31 249 35
rect 253 31 257 35
rect 271 31 275 35
rect 291 31 295 35
rect 303 31 307 35
rect 311 31 315 35
rect 329 31 333 35
rect 337 31 341 35
rect 355 31 359 35
rect 375 31 379 35
rect 387 31 391 35
rect 395 31 399 35
rect 406 31 410 35
rect 417 31 421 35
rect 425 31 429 35
rect 437 31 441 35
rect 445 31 449 35
rect 457 31 461 35
rect 475 31 479 35
rect 487 31 491 35
rect 495 31 499 35
rect 512 31 516 35
rect 523 31 527 35
rect 531 31 535 35
rect 543 31 547 35
rect 551 31 555 35
<< pdcontact >>
rect -32 269 -28 277
rect -24 269 -20 277
rect -6 269 -2 277
rect 2 269 6 277
rect 14 269 18 277
rect 26 269 30 277
rect 34 269 38 277
rect 52 269 56 277
rect 60 269 64 277
rect 78 269 82 277
rect 86 269 90 277
rect 98 269 102 277
rect 110 269 114 277
rect 118 269 122 277
rect 129 269 133 277
rect 148 269 152 277
rect 160 269 164 277
rect 168 269 172 277
rect 180 269 184 277
rect 188 269 194 277
rect 198 269 202 277
rect 210 269 214 277
rect 218 269 222 277
rect 245 269 249 277
rect 253 269 257 277
rect 271 269 275 277
rect 279 269 283 277
rect 291 269 295 277
rect 303 269 307 277
rect 311 269 315 277
rect 329 269 333 277
rect 337 269 341 277
rect 355 269 359 277
rect 363 269 367 277
rect 375 269 379 277
rect 387 269 391 277
rect 395 269 399 277
rect 406 269 410 277
rect 425 269 429 277
rect 437 269 441 277
rect 445 269 449 277
rect 457 269 461 277
rect 465 269 471 277
rect 475 269 479 277
rect 487 269 491 277
rect 495 269 499 277
rect 512 269 516 277
rect 531 269 535 277
rect 543 269 547 277
rect 551 269 555 277
rect -32 202 -28 210
rect -24 202 -20 210
rect -6 202 -2 210
rect 2 202 6 210
rect 14 202 18 210
rect 26 202 30 210
rect 34 202 38 210
rect 52 202 56 210
rect 60 202 64 210
rect 78 202 82 210
rect 86 202 90 210
rect 98 202 102 210
rect 110 202 114 210
rect 118 202 122 210
rect 129 202 133 210
rect 148 202 152 210
rect 160 202 164 210
rect 168 202 172 210
rect 180 202 184 210
rect 188 202 194 210
rect 198 202 202 210
rect 210 202 214 210
rect 218 202 222 210
rect 245 202 249 210
rect 253 202 257 210
rect 271 202 275 210
rect 279 202 283 210
rect 291 202 295 210
rect 303 202 307 210
rect 311 202 315 210
rect 329 202 333 210
rect 337 202 341 210
rect 355 202 359 210
rect 363 202 367 210
rect 375 202 379 210
rect 387 202 391 210
rect 395 202 399 210
rect 406 202 410 210
rect 425 202 429 210
rect 437 202 441 210
rect 445 202 449 210
rect 457 202 461 210
rect 465 202 471 210
rect 475 202 479 210
rect 487 202 491 210
rect 495 202 499 210
rect 512 202 516 210
rect 531 202 535 210
rect 543 202 547 210
rect 551 202 555 210
rect -32 135 -28 143
rect -24 135 -20 143
rect -6 135 -2 143
rect 2 135 6 143
rect 14 135 18 143
rect 26 135 30 143
rect 34 135 38 143
rect 52 135 56 143
rect 60 135 64 143
rect 78 135 82 143
rect 86 135 90 143
rect 98 135 102 143
rect 110 135 114 143
rect 118 135 122 143
rect 129 135 133 143
rect 148 135 152 143
rect 160 135 164 143
rect 168 135 172 143
rect 180 135 184 143
rect 188 135 194 143
rect 198 135 202 143
rect 210 135 214 143
rect 218 135 222 143
rect 245 135 249 143
rect 253 135 257 143
rect 271 135 275 143
rect 279 135 283 143
rect 291 135 295 143
rect 303 135 307 143
rect 311 135 315 143
rect 329 135 333 143
rect 337 135 341 143
rect 355 135 359 143
rect 363 135 367 143
rect 375 135 379 143
rect 387 135 391 143
rect 395 135 399 143
rect 406 135 410 143
rect 425 135 429 143
rect 437 135 441 143
rect 445 135 449 143
rect 457 135 461 143
rect 465 135 471 143
rect 475 135 479 143
rect 487 135 491 143
rect 495 135 499 143
rect 512 135 516 143
rect 531 135 535 143
rect 543 135 547 143
rect 551 135 555 143
rect -32 68 -28 76
rect -24 68 -20 76
rect -6 68 -2 76
rect 2 68 6 76
rect 14 68 18 76
rect 26 68 30 76
rect 34 68 38 76
rect 52 68 56 76
rect 60 68 64 76
rect 78 68 82 76
rect 86 68 90 76
rect 98 68 102 76
rect 110 68 114 76
rect 118 68 122 76
rect 129 68 133 76
rect 148 68 152 76
rect 160 68 164 76
rect 168 68 172 76
rect 180 68 184 76
rect 188 68 194 76
rect 198 68 202 76
rect 210 68 214 76
rect 218 68 222 76
rect 245 68 249 76
rect 253 68 257 76
rect 271 68 275 76
rect 279 68 283 76
rect 291 68 295 76
rect 303 68 307 76
rect 311 68 315 76
rect 329 68 333 76
rect 337 68 341 76
rect 355 68 359 76
rect 363 68 367 76
rect 375 68 379 76
rect 387 68 391 76
rect 395 68 399 76
rect 406 68 410 76
rect 425 68 429 76
rect 437 68 441 76
rect 445 68 449 76
rect 457 68 461 76
rect 465 68 471 76
rect 475 68 479 76
rect 487 68 491 76
rect 495 68 499 76
rect 512 68 516 76
rect 531 68 535 76
rect 543 68 547 76
rect 551 68 555 76
<< psubstratepcontact >>
rect -27 224 -18 228
rect -1 224 8 228
rect 31 224 40 228
rect 57 224 66 228
rect 83 224 92 228
rect 115 224 124 228
rect 165 224 174 228
rect 215 224 224 228
rect 250 224 259 228
rect 276 224 285 228
rect 308 224 317 228
rect 334 224 343 228
rect 360 224 369 228
rect 392 224 401 228
rect 442 224 451 228
rect 492 224 501 228
rect 548 224 557 228
rect -27 157 -18 161
rect -1 157 8 161
rect 31 157 40 161
rect 57 157 66 161
rect 83 157 92 161
rect 115 157 124 161
rect 165 157 174 161
rect 215 157 224 161
rect 250 157 259 161
rect 276 157 285 161
rect 308 157 317 161
rect 334 157 343 161
rect 360 157 369 161
rect 392 157 401 161
rect 442 157 451 161
rect 492 157 501 161
rect 548 157 557 161
rect -27 90 -18 94
rect -1 90 8 94
rect 31 90 40 94
rect 57 90 66 94
rect 83 90 92 94
rect 115 90 124 94
rect 165 90 174 94
rect 215 90 224 94
rect 250 90 259 94
rect 276 90 285 94
rect 308 90 317 94
rect 334 90 343 94
rect 360 90 369 94
rect 392 90 401 94
rect 442 90 451 94
rect 492 90 501 94
rect 548 90 557 94
rect -27 23 -18 27
rect -1 23 8 27
rect 31 23 40 27
rect 57 23 66 27
rect 83 23 92 27
rect 115 23 124 27
rect 165 23 174 27
rect 215 23 224 27
rect 250 23 259 27
rect 276 23 285 27
rect 308 23 317 27
rect 334 23 343 27
rect 360 23 369 27
rect 392 23 401 27
rect 442 23 451 27
rect 492 23 501 27
rect 548 23 557 27
<< nsubstratencontact >>
rect -27 281 -17 285
rect -1 281 9 285
rect 31 281 41 285
rect 57 281 67 285
rect 83 281 93 285
rect 115 281 125 285
rect 165 281 175 285
rect 215 281 225 285
rect 250 281 260 285
rect 276 281 286 285
rect 308 281 318 285
rect 334 281 344 285
rect 360 281 370 285
rect 392 281 402 285
rect 442 281 452 285
rect 492 281 502 285
rect 548 281 558 285
rect -27 214 -17 218
rect -1 214 9 218
rect 31 214 41 218
rect 57 214 67 218
rect 83 214 93 218
rect 115 214 125 218
rect 165 214 175 218
rect 215 214 225 218
rect 250 214 260 218
rect 276 214 286 218
rect 308 214 318 218
rect 334 214 344 218
rect 360 214 370 218
rect 392 214 402 218
rect 442 214 452 218
rect 492 214 502 218
rect 548 214 558 218
rect -27 147 -17 151
rect -1 147 9 151
rect 31 147 41 151
rect 57 147 67 151
rect 83 147 93 151
rect 115 147 125 151
rect 165 147 175 151
rect 215 147 225 151
rect 250 147 260 151
rect 276 147 286 151
rect 308 147 318 151
rect 334 147 344 151
rect 360 147 370 151
rect 392 147 402 151
rect 442 147 452 151
rect 492 147 502 151
rect 548 147 558 151
rect -27 80 -17 84
rect -1 80 9 84
rect 31 80 41 84
rect 57 80 67 84
rect 83 80 93 84
rect 115 80 125 84
rect 165 80 175 84
rect 215 80 225 84
rect 250 80 260 84
rect 276 80 286 84
rect 308 80 318 84
rect 334 80 344 84
rect 360 80 370 84
rect 392 80 402 84
rect 442 80 452 84
rect 492 80 502 84
rect 548 80 558 84
<< polysilicon >>
rect -27 277 -25 280
rect -1 277 1 280
rect 11 277 13 280
rect 31 277 33 280
rect 57 277 59 280
rect 83 277 85 280
rect 95 277 97 280
rect 115 277 117 280
rect 134 277 136 280
rect 145 277 147 280
rect 165 277 167 280
rect 185 277 187 280
rect 195 277 197 280
rect 215 277 217 280
rect 250 277 252 280
rect 276 277 278 280
rect 288 277 290 280
rect 308 277 310 280
rect 334 277 336 280
rect 360 277 362 280
rect 372 277 374 280
rect 392 277 394 280
rect 411 277 413 280
rect 422 277 424 280
rect 442 277 444 280
rect 462 277 464 280
rect 472 277 474 280
rect 492 277 494 280
rect 517 277 519 280
rect 528 277 530 280
rect 548 277 550 280
rect -27 236 -25 269
rect -1 236 1 269
rect 11 236 13 269
rect 31 236 33 269
rect 57 236 59 269
rect 83 236 85 269
rect 95 236 97 269
rect 115 236 117 269
rect 134 236 136 269
rect 145 236 147 269
rect 165 236 167 269
rect 185 236 187 269
rect 195 236 197 269
rect 215 236 217 269
rect 250 236 252 269
rect 276 236 278 269
rect 288 236 290 269
rect 308 236 310 269
rect 334 236 336 269
rect 360 236 362 269
rect 372 236 374 269
rect 392 236 394 269
rect 411 236 413 269
rect 422 236 424 269
rect 442 236 444 269
rect 462 236 464 269
rect 472 236 474 269
rect 492 236 494 269
rect 517 236 519 269
rect 528 236 530 269
rect 548 236 550 269
rect -27 229 -25 232
rect -1 229 1 232
rect 11 229 13 232
rect 31 229 33 232
rect 57 229 59 232
rect 83 229 85 232
rect 95 229 97 232
rect 115 229 117 232
rect 134 229 136 232
rect 145 229 147 232
rect 165 229 167 232
rect 185 229 187 232
rect 195 229 197 232
rect 215 229 217 232
rect 250 229 252 232
rect 276 229 278 232
rect 288 229 290 232
rect 308 229 310 232
rect 334 229 336 232
rect 360 229 362 232
rect 372 229 374 232
rect 392 229 394 232
rect 411 229 413 232
rect 422 229 424 232
rect 442 229 444 232
rect 462 229 464 232
rect 472 229 474 232
rect 492 229 494 232
rect 517 229 519 232
rect 528 229 530 232
rect 548 229 550 232
rect -27 210 -25 213
rect -1 210 1 213
rect 11 210 13 213
rect 31 210 33 213
rect 57 210 59 213
rect 83 210 85 213
rect 95 210 97 213
rect 115 210 117 213
rect 134 210 136 213
rect 145 210 147 213
rect 165 210 167 213
rect 185 210 187 213
rect 195 210 197 213
rect 215 210 217 213
rect 250 210 252 213
rect 276 210 278 213
rect 288 210 290 213
rect 308 210 310 213
rect 334 210 336 213
rect 360 210 362 213
rect 372 210 374 213
rect 392 210 394 213
rect 411 210 413 213
rect 422 210 424 213
rect 442 210 444 213
rect 462 210 464 213
rect 472 210 474 213
rect 492 210 494 213
rect 517 210 519 213
rect 528 210 530 213
rect 548 210 550 213
rect -27 169 -25 202
rect -1 169 1 202
rect 11 169 13 202
rect 31 169 33 202
rect 57 169 59 202
rect 83 169 85 202
rect 95 169 97 202
rect 115 169 117 202
rect 134 169 136 202
rect 145 169 147 202
rect 165 169 167 202
rect 185 169 187 202
rect 195 169 197 202
rect 215 169 217 202
rect 250 169 252 202
rect 276 169 278 202
rect 288 169 290 202
rect 308 169 310 202
rect 334 169 336 202
rect 360 169 362 202
rect 372 169 374 202
rect 392 169 394 202
rect 411 169 413 202
rect 422 169 424 202
rect 442 169 444 202
rect 462 169 464 202
rect 472 169 474 202
rect 492 169 494 202
rect 517 169 519 202
rect 528 169 530 202
rect 548 169 550 202
rect -27 162 -25 165
rect -1 162 1 165
rect 11 162 13 165
rect 31 162 33 165
rect 57 162 59 165
rect 83 162 85 165
rect 95 162 97 165
rect 115 162 117 165
rect 134 162 136 165
rect 145 162 147 165
rect 165 162 167 165
rect 185 162 187 165
rect 195 162 197 165
rect 215 162 217 165
rect 250 162 252 165
rect 276 162 278 165
rect 288 162 290 165
rect 308 162 310 165
rect 334 162 336 165
rect 360 162 362 165
rect 372 162 374 165
rect 392 162 394 165
rect 411 162 413 165
rect 422 162 424 165
rect 442 162 444 165
rect 462 162 464 165
rect 472 162 474 165
rect 492 162 494 165
rect 517 162 519 165
rect 528 162 530 165
rect 548 162 550 165
rect -27 143 -25 146
rect -1 143 1 146
rect 11 143 13 146
rect 31 143 33 146
rect 57 143 59 146
rect 83 143 85 146
rect 95 143 97 146
rect 115 143 117 146
rect 134 143 136 146
rect 145 143 147 146
rect 165 143 167 146
rect 185 143 187 146
rect 195 143 197 146
rect 215 143 217 146
rect 250 143 252 146
rect 276 143 278 146
rect 288 143 290 146
rect 308 143 310 146
rect 334 143 336 146
rect 360 143 362 146
rect 372 143 374 146
rect 392 143 394 146
rect 411 143 413 146
rect 422 143 424 146
rect 442 143 444 146
rect 462 143 464 146
rect 472 143 474 146
rect 492 143 494 146
rect 517 143 519 146
rect 528 143 530 146
rect 548 143 550 146
rect -27 102 -25 135
rect -1 102 1 135
rect 11 102 13 135
rect 31 102 33 135
rect 57 102 59 135
rect 83 102 85 135
rect 95 102 97 135
rect 115 102 117 135
rect 134 102 136 135
rect 145 102 147 135
rect 165 102 167 135
rect 185 102 187 135
rect 195 102 197 135
rect 215 102 217 135
rect 250 102 252 135
rect 276 102 278 135
rect 288 102 290 135
rect 308 102 310 135
rect 334 102 336 135
rect 360 102 362 135
rect 372 102 374 135
rect 392 102 394 135
rect 411 102 413 135
rect 422 102 424 135
rect 442 102 444 135
rect 462 102 464 135
rect 472 102 474 135
rect 492 102 494 135
rect 517 102 519 135
rect 528 102 530 135
rect 548 102 550 135
rect -27 95 -25 98
rect -1 95 1 98
rect 11 95 13 98
rect 31 95 33 98
rect 57 95 59 98
rect 83 95 85 98
rect 95 95 97 98
rect 115 95 117 98
rect 134 95 136 98
rect 145 95 147 98
rect 165 95 167 98
rect 185 95 187 98
rect 195 95 197 98
rect 215 95 217 98
rect 250 95 252 98
rect 276 95 278 98
rect 288 95 290 98
rect 308 95 310 98
rect 334 95 336 98
rect 360 95 362 98
rect 372 95 374 98
rect 392 95 394 98
rect 411 95 413 98
rect 422 95 424 98
rect 442 95 444 98
rect 462 95 464 98
rect 472 95 474 98
rect 492 95 494 98
rect 517 95 519 98
rect 528 95 530 98
rect 548 95 550 98
rect -27 76 -25 79
rect -1 76 1 79
rect 11 76 13 79
rect 31 76 33 79
rect 57 76 59 79
rect 83 76 85 79
rect 95 76 97 79
rect 115 76 117 79
rect 134 76 136 79
rect 145 76 147 79
rect 165 76 167 79
rect 185 76 187 79
rect 195 76 197 79
rect 215 76 217 79
rect 250 76 252 79
rect 276 76 278 79
rect 288 76 290 79
rect 308 76 310 79
rect 334 76 336 79
rect 360 76 362 79
rect 372 76 374 79
rect 392 76 394 79
rect 411 76 413 79
rect 422 76 424 79
rect 442 76 444 79
rect 462 76 464 79
rect 472 76 474 79
rect 492 76 494 79
rect 517 76 519 79
rect 528 76 530 79
rect 548 76 550 79
rect -27 35 -25 68
rect -1 35 1 68
rect 11 35 13 68
rect 31 35 33 68
rect 57 35 59 68
rect 83 35 85 68
rect 95 35 97 68
rect 115 35 117 68
rect 134 35 136 68
rect 145 35 147 68
rect 165 35 167 68
rect 185 35 187 68
rect 195 35 197 68
rect 215 35 217 68
rect 250 35 252 68
rect 276 35 278 68
rect 288 35 290 68
rect 308 35 310 68
rect 334 35 336 68
rect 360 35 362 68
rect 372 35 374 68
rect 392 35 394 68
rect 411 35 413 68
rect 422 35 424 68
rect 442 35 444 68
rect 462 35 464 68
rect 472 35 474 68
rect 492 35 494 68
rect 517 35 519 68
rect 528 35 530 68
rect 548 35 550 68
rect -27 28 -25 31
rect -1 28 1 31
rect 11 28 13 31
rect 31 28 33 31
rect 57 28 59 31
rect 83 28 85 31
rect 95 28 97 31
rect 115 28 117 31
rect 134 28 136 31
rect 145 28 147 31
rect 165 28 167 31
rect 185 28 187 31
rect 195 28 197 31
rect 215 28 217 31
rect 250 28 252 31
rect 276 28 278 31
rect 288 28 290 31
rect 308 28 310 31
rect 334 28 336 31
rect 360 28 362 31
rect 372 28 374 31
rect 392 28 394 31
rect 411 28 413 31
rect 422 28 424 31
rect 442 28 444 31
rect 462 28 464 31
rect 472 28 474 31
rect 492 28 494 31
rect 517 28 519 31
rect 528 28 530 31
rect 548 28 550 31
<< polycontact >>
rect -31 261 -27 265
rect -5 261 -1 265
rect 7 254 11 258
rect 27 261 31 265
rect 53 261 57 265
rect 79 261 83 265
rect 91 237 95 241
rect 111 261 115 265
rect 130 246 134 250
rect 141 262 145 266
rect 161 261 165 265
rect 181 261 185 265
rect 191 239 195 243
rect 210 261 215 266
rect 246 261 250 265
rect 272 261 276 265
rect 284 254 288 258
rect 304 261 308 265
rect 330 261 334 265
rect 356 261 360 265
rect 368 237 372 241
rect 388 261 392 265
rect 407 246 411 250
rect 418 262 422 266
rect 438 261 442 265
rect 458 261 462 265
rect 468 239 472 243
rect 487 261 492 266
rect 513 246 517 250
rect 524 262 528 266
rect 544 261 548 265
rect -31 194 -27 198
rect -5 194 -1 198
rect 7 187 11 191
rect 27 194 31 198
rect 53 194 57 198
rect 79 194 83 198
rect 91 170 95 174
rect 111 194 115 198
rect 130 179 134 183
rect 141 195 145 199
rect 161 194 165 198
rect 181 194 185 198
rect 191 172 195 176
rect 210 194 215 199
rect 246 194 250 198
rect 272 194 276 198
rect 284 187 288 191
rect 304 194 308 198
rect 330 194 334 198
rect 356 194 360 198
rect 368 170 372 174
rect 388 194 392 198
rect 407 179 411 183
rect 418 195 422 199
rect 438 194 442 198
rect 458 194 462 198
rect 468 172 472 176
rect 487 194 492 199
rect 513 179 517 183
rect 524 195 528 199
rect 544 194 548 198
rect -31 127 -27 131
rect -5 127 -1 131
rect 7 120 11 124
rect 27 127 31 131
rect 53 127 57 131
rect 79 127 83 131
rect 91 103 95 107
rect 111 127 115 131
rect 130 112 134 116
rect 141 128 145 132
rect 161 127 165 131
rect 181 127 185 131
rect 191 105 195 109
rect 210 127 215 132
rect 246 127 250 131
rect 272 127 276 131
rect 284 120 288 124
rect 304 127 308 131
rect 330 127 334 131
rect 356 127 360 131
rect 368 103 372 107
rect 388 127 392 131
rect 407 112 411 116
rect 418 128 422 132
rect 438 127 442 131
rect 458 127 462 131
rect 468 105 472 109
rect 487 127 492 132
rect 513 112 517 116
rect 524 128 528 132
rect 544 127 548 131
rect -31 60 -27 64
rect -5 60 -1 64
rect 7 53 11 57
rect 27 60 31 64
rect 53 60 57 64
rect 79 60 83 64
rect 91 36 95 40
rect 111 60 115 64
rect 130 45 134 49
rect 141 61 145 65
rect 161 60 165 64
rect 181 60 185 64
rect 191 38 195 42
rect 210 60 215 65
rect 246 60 250 64
rect 272 60 276 64
rect 284 53 288 57
rect 304 60 308 64
rect 330 60 334 64
rect 356 60 360 64
rect 368 36 372 40
rect 388 60 392 64
rect 407 45 411 49
rect 418 61 422 65
rect 438 60 442 64
rect 458 60 462 64
rect 468 38 472 42
rect 487 60 492 65
rect 513 45 517 49
rect 524 61 528 65
rect 544 60 548 64
<< metal1 >>
rect -36 285 569 286
rect -36 281 -27 285
rect -17 281 -1 285
rect 9 281 31 285
rect 41 281 57 285
rect 67 281 83 285
rect 93 281 115 285
rect 125 281 165 285
rect 175 281 215 285
rect 225 281 250 285
rect 260 281 276 285
rect 286 281 308 285
rect 318 281 334 285
rect 344 281 360 285
rect 370 281 392 285
rect 402 281 442 285
rect 452 281 492 285
rect 502 281 548 285
rect 558 281 569 285
rect -32 277 -28 281
rect -6 277 -2 281
rect 14 277 18 281
rect 26 277 30 281
rect 52 277 56 281
rect 78 277 82 281
rect 98 277 102 281
rect 110 277 114 281
rect 129 277 133 281
rect 160 277 164 281
rect 180 277 184 281
rect 198 277 202 281
rect 210 277 214 281
rect 245 277 249 281
rect 271 277 275 281
rect 291 277 295 281
rect 303 277 307 281
rect 329 277 333 281
rect 355 277 359 281
rect 375 277 379 281
rect 387 277 391 281
rect 406 277 410 281
rect 437 277 441 281
rect 457 277 461 281
rect 475 277 479 281
rect 487 277 491 281
rect 512 277 516 281
rect 543 277 547 281
rect -24 265 -20 269
rect 2 265 6 269
rect -38 261 -36 265
rect -24 261 -5 265
rect 2 261 27 265
rect -24 236 -20 261
rect -8 254 2 258
rect 14 236 18 261
rect 34 250 38 269
rect 60 265 64 269
rect 86 265 90 269
rect 118 266 122 269
rect 60 261 79 265
rect 86 261 111 265
rect 118 262 141 266
rect 148 265 152 269
rect 34 236 38 245
rect 60 236 64 261
rect 98 236 102 261
rect 118 236 122 262
rect 148 261 161 265
rect 148 259 152 261
rect 140 255 152 259
rect 140 236 144 255
rect 168 236 172 269
rect 188 266 194 269
rect 188 261 210 266
rect 198 236 203 261
rect 218 236 222 269
rect 253 265 257 269
rect 279 265 283 269
rect 239 261 241 265
rect 253 261 272 265
rect 279 261 304 265
rect 253 236 257 261
rect 269 254 279 258
rect 291 236 295 261
rect 311 250 315 269
rect 337 265 341 269
rect 363 265 367 269
rect 395 266 399 269
rect 337 261 356 265
rect 363 261 388 265
rect 395 262 418 266
rect 425 265 429 269
rect 311 236 315 245
rect 337 236 341 261
rect 375 236 379 261
rect 395 236 399 262
rect 425 261 438 265
rect 425 259 429 261
rect 417 255 429 259
rect 445 257 449 269
rect 465 266 471 269
rect 495 266 499 269
rect 465 261 487 266
rect 495 262 524 266
rect 531 265 535 269
rect 417 236 421 255
rect 445 253 454 257
rect 445 236 449 253
rect 475 236 480 261
rect 495 236 499 262
rect 531 261 544 265
rect 531 259 535 261
rect 523 255 535 259
rect 523 236 527 255
rect 551 236 555 269
rect -32 228 -28 232
rect -6 228 -2 232
rect 26 228 30 232
rect 52 228 56 232
rect 78 228 82 232
rect 110 228 114 232
rect 129 228 133 232
rect 148 228 152 232
rect 202 232 203 236
rect 160 228 164 232
rect 180 228 184 232
rect 210 228 214 232
rect 245 228 249 232
rect 271 228 275 232
rect 303 228 307 232
rect 329 228 333 232
rect 355 228 359 232
rect 387 228 391 232
rect 406 228 410 232
rect 425 228 429 232
rect 479 232 480 236
rect 437 228 441 232
rect 457 228 461 232
rect 487 228 491 232
rect 512 228 516 232
rect 531 228 535 232
rect 543 228 547 232
rect -46 224 -27 228
rect -18 224 -1 228
rect 8 224 31 228
rect 40 224 57 228
rect 66 224 83 228
rect 92 224 115 228
rect 124 224 165 228
rect 174 224 215 228
rect 224 224 250 228
rect 259 224 276 228
rect 285 224 308 228
rect 317 224 334 228
rect 343 224 360 228
rect 369 224 392 228
rect 401 224 442 228
rect 451 224 492 228
rect 501 224 548 228
rect 557 224 562 228
rect -46 223 562 224
rect -46 161 -42 223
rect 565 219 569 281
rect -36 218 569 219
rect -36 214 -27 218
rect -17 214 -1 218
rect 9 214 31 218
rect 41 214 57 218
rect 67 214 83 218
rect 93 214 115 218
rect 125 214 165 218
rect 175 214 215 218
rect 225 214 250 218
rect 260 214 276 218
rect 286 214 308 218
rect 318 214 334 218
rect 344 214 360 218
rect 370 214 392 218
rect 402 214 442 218
rect 452 214 492 218
rect 502 214 548 218
rect 558 214 569 218
rect -32 210 -28 214
rect -6 210 -2 214
rect 14 210 18 214
rect 26 210 30 214
rect 52 210 56 214
rect 78 210 82 214
rect 98 210 102 214
rect 110 210 114 214
rect 129 210 133 214
rect 160 210 164 214
rect 180 210 184 214
rect 198 210 202 214
rect 210 210 214 214
rect 245 210 249 214
rect 271 210 275 214
rect 291 210 295 214
rect 303 210 307 214
rect 329 210 333 214
rect 355 210 359 214
rect 375 210 379 214
rect 387 210 391 214
rect 406 210 410 214
rect 437 210 441 214
rect 457 210 461 214
rect 475 210 479 214
rect 487 210 491 214
rect 512 210 516 214
rect 543 210 547 214
rect -24 198 -20 202
rect 2 198 6 202
rect -38 194 -36 198
rect -24 194 -5 198
rect 2 194 27 198
rect -24 169 -20 194
rect -8 187 2 191
rect 14 169 18 194
rect 34 183 38 202
rect 60 198 64 202
rect 86 198 90 202
rect 118 199 122 202
rect 60 194 79 198
rect 86 194 111 198
rect 118 195 141 199
rect 148 198 152 202
rect 34 169 38 178
rect 60 169 64 194
rect 98 169 102 194
rect 118 169 122 195
rect 148 194 161 198
rect 148 192 152 194
rect 140 188 152 192
rect 140 169 144 188
rect 168 169 172 202
rect 188 199 194 202
rect 188 194 210 199
rect 198 169 203 194
rect 218 169 222 202
rect 253 198 257 202
rect 279 198 283 202
rect 239 194 241 198
rect 253 194 272 198
rect 279 194 304 198
rect 253 169 257 194
rect 273 187 279 191
rect 291 169 295 194
rect 311 183 315 202
rect 337 198 341 202
rect 363 198 367 202
rect 395 199 399 202
rect 337 194 356 198
rect 363 194 388 198
rect 395 195 418 199
rect 425 198 429 202
rect 311 169 315 178
rect 337 169 341 194
rect 375 169 379 194
rect 395 169 399 195
rect 425 194 438 198
rect 425 192 429 194
rect 417 188 429 192
rect 445 190 449 202
rect 465 199 471 202
rect 495 199 499 202
rect 465 194 487 199
rect 495 195 524 199
rect 531 198 535 202
rect 417 169 421 188
rect 445 186 454 190
rect 445 169 449 186
rect 475 169 480 194
rect 495 169 499 195
rect 531 194 544 198
rect 531 192 535 194
rect 523 188 535 192
rect 523 169 527 188
rect 551 169 555 202
rect -32 161 -28 165
rect -6 161 -2 165
rect 26 161 30 165
rect 52 161 56 165
rect 78 161 82 165
rect 110 161 114 165
rect 129 161 133 165
rect 148 161 152 165
rect 202 165 203 169
rect 160 161 164 165
rect 180 161 184 165
rect 210 161 214 165
rect 245 161 249 165
rect 271 161 275 165
rect 303 161 307 165
rect 329 161 333 165
rect 355 161 359 165
rect 387 161 391 165
rect 406 161 410 165
rect 425 161 429 165
rect 479 165 480 169
rect 437 161 441 165
rect 457 161 461 165
rect 487 161 491 165
rect 512 161 516 165
rect 531 161 535 165
rect 543 161 547 165
rect -46 157 -27 161
rect -18 157 -1 161
rect 8 157 31 161
rect 40 157 57 161
rect 66 157 83 161
rect 92 157 115 161
rect 124 157 165 161
rect 174 157 215 161
rect 224 157 250 161
rect 259 157 276 161
rect 285 157 308 161
rect 317 157 334 161
rect 343 157 360 161
rect 369 157 392 161
rect 401 157 442 161
rect 451 157 492 161
rect 501 157 548 161
rect 557 157 562 161
rect -46 156 562 157
rect -46 94 -42 156
rect 565 152 569 214
rect -36 151 569 152
rect -36 147 -27 151
rect -17 147 -1 151
rect 9 147 31 151
rect 41 147 57 151
rect 67 147 83 151
rect 93 147 115 151
rect 125 147 165 151
rect 175 147 215 151
rect 225 147 250 151
rect 260 147 276 151
rect 286 147 308 151
rect 318 147 334 151
rect 344 147 360 151
rect 370 147 392 151
rect 402 147 442 151
rect 452 147 492 151
rect 502 147 548 151
rect 558 147 569 151
rect -32 143 -28 147
rect -6 143 -2 147
rect 14 143 18 147
rect 26 143 30 147
rect 52 143 56 147
rect 78 143 82 147
rect 98 143 102 147
rect 110 143 114 147
rect 129 143 133 147
rect 160 143 164 147
rect 180 143 184 147
rect 198 143 202 147
rect 210 143 214 147
rect 245 143 249 147
rect 271 143 275 147
rect 291 143 295 147
rect 303 143 307 147
rect 329 143 333 147
rect 355 143 359 147
rect 375 143 379 147
rect 387 143 391 147
rect 406 143 410 147
rect 437 143 441 147
rect 457 143 461 147
rect 475 143 479 147
rect 487 143 491 147
rect 512 143 516 147
rect 543 143 547 147
rect -24 131 -20 135
rect 2 131 6 135
rect -39 127 -36 131
rect -24 127 -5 131
rect 2 127 27 131
rect -24 102 -20 127
rect -8 120 2 124
rect 14 102 18 127
rect 34 116 38 135
rect 60 131 64 135
rect 86 131 90 135
rect 118 132 122 135
rect 60 127 79 131
rect 86 127 111 131
rect 118 128 141 132
rect 148 131 152 135
rect 34 102 38 111
rect 60 102 64 127
rect 98 102 102 127
rect 118 102 122 128
rect 148 127 161 131
rect 148 125 152 127
rect 140 121 152 125
rect 140 102 144 121
rect 168 102 172 135
rect 188 132 194 135
rect 188 127 210 132
rect 198 102 203 127
rect 218 102 222 135
rect 253 131 257 135
rect 279 131 283 135
rect 239 127 241 131
rect 253 127 272 131
rect 279 127 304 131
rect 253 102 257 127
rect 272 120 279 124
rect 291 102 295 127
rect 311 116 315 135
rect 337 131 341 135
rect 363 131 367 135
rect 395 132 399 135
rect 337 127 356 131
rect 363 127 388 131
rect 395 128 418 132
rect 425 131 429 135
rect 311 102 315 111
rect 337 102 341 127
rect 375 102 379 127
rect 395 102 399 128
rect 425 127 438 131
rect 425 125 429 127
rect 417 121 429 125
rect 445 123 449 135
rect 465 132 471 135
rect 495 132 499 135
rect 465 127 487 132
rect 495 128 524 132
rect 531 131 535 135
rect 417 102 421 121
rect 445 119 454 123
rect 445 102 449 119
rect 475 102 480 127
rect 495 102 499 128
rect 531 127 544 131
rect 531 125 535 127
rect 523 121 535 125
rect 523 102 527 121
rect 551 102 555 135
rect -32 94 -28 98
rect -6 94 -2 98
rect 26 94 30 98
rect 52 94 56 98
rect 78 94 82 98
rect 110 94 114 98
rect 129 94 133 98
rect 148 94 152 98
rect 202 98 203 102
rect 160 94 164 98
rect 180 94 184 98
rect 210 94 214 98
rect 245 94 249 98
rect 271 94 275 98
rect 303 94 307 98
rect 329 94 333 98
rect 355 94 359 98
rect 387 94 391 98
rect 406 94 410 98
rect 425 94 429 98
rect 479 98 480 102
rect 437 94 441 98
rect 457 94 461 98
rect 487 94 491 98
rect 512 94 516 98
rect 531 94 535 98
rect 543 94 547 98
rect -46 90 -27 94
rect -18 90 -1 94
rect 8 90 31 94
rect 40 90 57 94
rect 66 90 83 94
rect 92 90 115 94
rect 124 90 165 94
rect 174 90 215 94
rect 224 90 250 94
rect 259 90 276 94
rect 285 90 308 94
rect 317 90 334 94
rect 343 90 360 94
rect 369 90 392 94
rect 401 90 442 94
rect 451 90 492 94
rect 501 90 548 94
rect 557 90 562 94
rect -46 89 562 90
rect -46 27 -42 89
rect 565 85 569 147
rect -36 84 569 85
rect -36 80 -27 84
rect -17 80 -1 84
rect 9 80 31 84
rect 41 80 57 84
rect 67 80 83 84
rect 93 80 115 84
rect 125 80 165 84
rect 175 80 215 84
rect 225 80 250 84
rect 260 80 276 84
rect 286 80 308 84
rect 318 80 334 84
rect 344 80 360 84
rect 370 80 392 84
rect 402 80 442 84
rect 452 80 492 84
rect 502 80 548 84
rect 558 80 569 84
rect -32 76 -28 80
rect -6 76 -2 80
rect 14 76 18 80
rect 26 76 30 80
rect 52 76 56 80
rect 78 76 82 80
rect 98 76 102 80
rect 110 76 114 80
rect 129 76 133 80
rect 160 76 164 80
rect 180 76 184 80
rect 198 76 202 80
rect 210 76 214 80
rect 245 76 249 80
rect 271 76 275 80
rect 291 76 295 80
rect 303 76 307 80
rect 329 76 333 80
rect 355 76 359 80
rect 375 76 379 80
rect 387 76 391 80
rect 406 76 410 80
rect 437 76 441 80
rect 457 76 461 80
rect 475 76 479 80
rect 487 76 491 80
rect 512 76 516 80
rect 543 76 547 80
rect -24 64 -20 68
rect 2 64 6 68
rect -39 60 -36 64
rect -24 60 -5 64
rect 2 60 27 64
rect -24 35 -20 60
rect -8 53 2 57
rect 14 35 18 60
rect 34 49 38 68
rect 60 64 64 68
rect 86 64 90 68
rect 118 65 122 68
rect 60 60 79 64
rect 86 60 111 64
rect 118 61 141 65
rect 148 64 152 68
rect 34 35 38 44
rect 60 35 64 60
rect 98 35 102 60
rect 118 35 122 61
rect 148 60 161 64
rect 148 58 152 60
rect 140 54 152 58
rect 140 35 144 54
rect 168 35 172 68
rect 188 65 194 68
rect 188 60 210 65
rect 198 35 203 60
rect 218 35 222 68
rect 253 64 257 68
rect 279 64 283 68
rect 239 60 241 64
rect 253 60 272 64
rect 279 60 304 64
rect 253 35 257 60
rect 272 53 279 57
rect 291 35 295 60
rect 311 49 315 68
rect 337 64 341 68
rect 363 64 367 68
rect 395 65 399 68
rect 337 60 356 64
rect 363 60 388 64
rect 395 61 418 65
rect 425 64 429 68
rect 311 35 315 44
rect 337 35 341 60
rect 375 35 379 60
rect 395 35 399 61
rect 425 60 438 64
rect 425 58 429 60
rect 417 54 429 58
rect 445 56 449 68
rect 465 65 471 68
rect 495 65 499 68
rect 465 60 487 65
rect 495 61 524 65
rect 531 64 535 68
rect 417 35 421 54
rect 445 52 454 56
rect 445 35 449 52
rect 475 35 480 60
rect 495 35 499 61
rect 531 60 544 64
rect 531 58 535 60
rect 523 54 535 58
rect 551 54 555 68
rect 523 35 527 54
rect 551 50 558 54
rect 551 35 555 50
rect -32 27 -28 31
rect -6 27 -2 31
rect 26 27 30 31
rect 52 27 56 31
rect 78 27 82 31
rect 110 27 114 31
rect 129 27 133 31
rect 148 27 152 31
rect 202 31 203 35
rect 160 27 164 31
rect 180 27 184 31
rect 210 27 214 31
rect 245 27 249 31
rect 271 27 275 31
rect 303 27 307 31
rect 329 27 333 31
rect 355 27 359 31
rect 387 27 391 31
rect 406 27 410 31
rect 425 27 429 31
rect 479 31 480 35
rect 437 27 441 31
rect 457 27 461 31
rect 487 27 491 31
rect 512 27 516 31
rect 531 27 535 31
rect 543 27 547 31
rect -46 23 -27 27
rect -18 23 -1 27
rect 8 23 31 27
rect 40 23 57 27
rect 66 23 83 27
rect 92 23 115 27
rect 124 23 165 27
rect 174 23 215 27
rect 224 23 250 27
rect 259 23 276 27
rect 285 23 308 27
rect 317 23 334 27
rect 343 23 360 27
rect 369 23 392 27
rect 401 23 442 27
rect 451 23 492 27
rect 501 23 548 27
rect -46 22 557 23
<< m2contact >>
rect -36 260 -31 265
rect 2 253 7 258
rect 48 260 53 265
rect 34 245 39 250
rect 86 237 91 242
rect 125 245 130 250
rect 176 260 181 265
rect 172 251 177 256
rect 186 239 191 244
rect 241 260 246 265
rect 222 237 227 242
rect 279 253 284 258
rect 325 260 330 265
rect 311 245 316 250
rect 363 237 368 242
rect 453 260 458 265
rect 402 245 407 250
rect 463 239 468 244
rect 508 245 513 250
rect 555 251 560 256
rect -36 193 -31 198
rect 2 186 7 191
rect 48 193 53 198
rect 34 178 39 183
rect 86 170 91 175
rect 125 178 130 183
rect 176 193 181 198
rect 172 184 177 189
rect 186 172 191 177
rect 241 193 246 198
rect 222 170 227 175
rect 279 186 284 191
rect 325 193 330 198
rect 311 178 316 183
rect 363 170 368 175
rect 453 193 458 198
rect 402 178 407 183
rect 463 172 468 177
rect 508 178 513 183
rect 555 184 560 189
rect -36 126 -31 131
rect 2 119 7 124
rect 48 126 53 131
rect 34 111 39 116
rect 86 103 91 108
rect 125 111 130 116
rect 176 126 181 131
rect 172 117 177 122
rect 186 105 191 110
rect 241 126 246 131
rect 222 103 227 108
rect 279 119 284 124
rect 325 126 330 131
rect 311 111 316 116
rect 363 103 368 108
rect 453 126 458 131
rect 402 111 407 116
rect 463 105 468 110
rect 508 111 513 116
rect 555 117 560 122
rect -36 59 -31 64
rect 2 52 7 57
rect 48 59 53 64
rect 34 44 39 49
rect 86 36 91 41
rect 125 44 130 49
rect 176 59 181 64
rect 172 50 177 55
rect 186 38 191 43
rect 241 59 246 64
rect 222 36 227 41
rect 279 52 284 57
rect 325 59 330 64
rect 311 44 316 49
rect 363 36 368 41
rect 453 59 458 64
rect 402 44 407 49
rect 463 38 468 43
rect 508 44 513 49
<< metal2 >>
rect -36 241 -31 260
rect 48 258 53 260
rect 74 261 176 265
rect 74 258 78 261
rect 7 254 78 258
rect 241 255 246 260
rect 325 258 330 260
rect 351 261 453 265
rect 351 258 355 261
rect 177 251 246 255
rect 284 254 355 258
rect 39 246 125 250
rect 130 246 134 250
rect -36 237 86 241
rect 175 241 186 243
rect 91 239 186 241
rect 91 237 180 239
rect 227 228 231 242
rect 241 241 246 251
rect 316 246 402 250
rect 407 246 411 250
rect 241 237 363 241
rect 452 241 463 243
rect 368 239 463 241
rect 368 237 457 239
rect 504 228 508 250
rect 227 224 508 228
rect 555 218 559 251
rect 279 214 559 218
rect -36 174 -31 193
rect 48 191 53 193
rect 74 194 176 198
rect 74 191 78 194
rect 7 187 78 191
rect 241 188 246 193
rect 177 184 246 188
rect 279 191 284 214
rect 325 191 330 193
rect 351 194 453 198
rect 351 191 355 194
rect 284 187 355 191
rect 39 179 125 183
rect 130 179 134 183
rect -36 170 86 174
rect 175 174 186 176
rect 91 172 186 174
rect 91 170 180 172
rect 227 161 231 175
rect 241 174 246 184
rect 316 179 402 183
rect 407 179 411 183
rect 241 170 363 174
rect 452 174 463 176
rect 368 172 463 174
rect 368 170 457 172
rect 504 161 508 183
rect 227 157 508 161
rect 555 151 559 184
rect 279 147 559 151
rect -36 107 -31 126
rect 48 124 53 126
rect 74 127 176 131
rect 74 124 78 127
rect 7 120 78 124
rect 241 121 246 126
rect 177 117 246 121
rect 279 124 284 147
rect 325 124 330 126
rect 351 127 453 131
rect 351 124 355 127
rect 284 120 355 124
rect 39 112 125 116
rect 130 112 134 116
rect -36 103 86 107
rect 175 107 186 109
rect 91 105 186 107
rect 91 103 180 105
rect 227 94 231 108
rect 241 107 246 117
rect 316 112 402 116
rect 407 112 411 116
rect 241 103 363 107
rect 452 107 463 109
rect 368 105 463 107
rect 368 103 457 105
rect 504 94 508 116
rect 227 90 508 94
rect 555 84 559 117
rect 279 80 559 84
rect -36 40 -31 59
rect 48 57 53 59
rect 74 60 176 64
rect 74 57 78 60
rect 7 53 78 57
rect 241 54 246 59
rect 177 50 246 54
rect 279 57 284 80
rect 325 57 330 59
rect 351 60 453 64
rect 351 57 355 60
rect 284 53 355 57
rect 39 45 125 49
rect 130 45 134 49
rect -36 36 86 40
rect 175 40 186 42
rect 91 38 186 40
rect 91 36 180 38
rect 227 27 231 41
rect 241 40 246 50
rect 316 45 402 49
rect 407 45 411 49
rect 241 36 363 40
rect 452 40 463 42
rect 368 38 463 40
rect 368 36 457 38
rect 504 27 508 49
rect 227 23 508 27
<< labels >>
rlabel metal1 -9 83 -9 83 4 Vdd
rlabel metal1 -10 25 -10 25 2 Gnd
rlabel metal1 268 83 268 83 4 Vdd
rlabel metal1 267 25 267 25 2 Gnd
rlabel metal1 -9 150 -9 150 4 Vdd
rlabel metal1 -10 92 -10 92 2 Gnd
rlabel metal1 268 150 268 150 4 Vdd
rlabel metal1 267 92 267 92 2 Gnd
rlabel metal1 -9 217 -9 217 4 Vdd
rlabel metal1 -10 159 -10 159 2 Gnd
rlabel metal1 268 217 268 217 4 Vdd
rlabel metal1 267 159 267 159 2 Gnd
rlabel metal1 -9 284 -9 284 4 Vdd
rlabel metal1 -10 226 -10 226 2 Gnd
rlabel metal1 268 284 268 284 4 Vdd
rlabel metal1 267 226 267 226 2 Gnd
rlabel metal1 271 255 271 255 1 Cin
rlabel m2contact -34 262 -34 262 3 A0
rlabel metal1 -6 255 -6 255 1 B0
rlabel m2contact -34 195 -34 195 3 A1
rlabel metal1 -6 189 -6 189 1 B1
rlabel m2contact -35 128 -35 128 3 A2
rlabel metal1 -5 121 -5 121 1 B2
rlabel metal1 -6 54 -6 54 1 B3
rlabel m2contact -33 61 -33 61 1 A3
rlabel metal1 452 255 452 255 1 S0
rlabel metal1 450 187 450 187 1 S1
rlabel metal1 451 121 451 121 1 S2
rlabel metal1 451 54 451 54 1 S3
rlabel metal1 556 52 556 52 1 Cout
<< end >>
