magic
tech scmos
timestamp 1699467758
<< nwell >>
rect -10 3 18 27
<< ntransistor >>
rect 2 -15 4 -11
<< ptransistor >>
rect 2 9 4 13
<< ndiffusion >>
rect 1 -15 2 -11
rect 4 -15 5 -11
rect 9 -15 10 -11
<< pdiffusion >>
rect 1 9 2 13
rect 4 9 5 13
rect 9 9 10 13
<< ndcontact >>
rect -3 -15 1 -11
rect 5 -15 9 -11
<< pdcontact >>
rect -3 9 1 13
rect 5 9 9 13
<< psubstratepcontact >>
rect -3 -24 1 -20
<< nsubstratencontact >>
rect -3 20 1 24
<< polysilicon >>
rect 2 13 4 16
rect 2 -2 4 9
rect 1 -6 4 -2
rect 2 -11 4 -6
rect 2 -18 4 -15
<< polycontact >>
rect -3 -6 1 -2
<< metal1 >>
rect -7 20 -3 24
rect 1 20 12 24
rect -3 13 1 20
rect 5 -2 9 9
rect -10 -6 -3 -2
rect 5 -6 14 -2
rect 5 -11 9 -6
rect -3 -20 1 -15
rect 1 -24 12 -20
<< labels >>
rlabel metal1 -10 -6 -10 -2 3 in
rlabel metal1 14 -6 14 -2 7 out
rlabel metal1 5 22 5 22 5 vdd!
rlabel metal1 5 -22 5 -22 1 gnd!
<< end >>
