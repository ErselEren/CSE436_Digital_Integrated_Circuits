* SPICE3 file created from test1.ext - technology: scmos

.option scale=0.12u

M1000 out in vdd vdd PMOS w=8 l=2
+  ad=64p pd=32u as=40p ps=26u
M1001 out in gnd Gnd NMOS w=4 l=2
+  ad=32p pd=24u as=20p ps=18u

.include tsmc_cmos025

Vs Vdd Gnd 2.5V
Vp in Gnd PULSE(0 2.5 2n 0.1n 0.1n 4n 10n)

.TRAN 1n 60n
.OPTIONS
