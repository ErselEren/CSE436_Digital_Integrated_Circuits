magic
tech scmos
timestamp 1699388788
<< nwell >>
rect -10 3 18 30
<< ntransistor >>
rect 2 -15 4 -11
<< ptransistor >>
rect 2 9 4 17
<< ndiffusion >>
rect 1 -15 2 -11
rect 4 -15 5 -11
rect 9 -15 12 -11
<< pdiffusion >>
rect 1 9 2 17
rect 4 9 5 17
rect 9 9 12 17
<< ndcontact >>
rect -3 -15 1 -11
rect 5 -15 9 -11
<< pdcontact >>
rect -3 9 1 17
rect 5 9 9 17
<< psubstratepcontact >>
rect -3 -24 1 -20
<< nsubstratencontact >>
rect -3 23 1 27
<< polysilicon >>
rect 2 17 4 20
rect 2 2 4 9
rect 0 0 4 2
rect 0 -2 2 0
rect 1 -6 2 -2
rect 0 -7 2 -6
rect 0 -9 4 -7
rect 2 -11 4 -9
rect 2 -18 4 -15
<< polycontact >>
rect -3 -6 1 -2
<< metal1 >>
rect -7 23 -3 27
rect 1 23 12 27
rect -3 17 1 23
rect 5 -2 9 9
rect -9 -6 -3 -2
rect 5 -6 14 -2
rect 5 -11 9 -6
rect -3 -20 1 -15
rect 1 -24 12 -20
<< labels >>
rlabel metal1 -9 -6 -9 -2 3 in
rlabel metal1 14 -6 14 -2 7 out
rlabel metal1 4 -22 4 -22 1 gnd!
rlabel metal1 3 25 3 25 5 vdd!
<< end >>
